VerbForm=Stem
